import uvm_pkg::*;
