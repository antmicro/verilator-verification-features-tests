/*
:name: easyUVM
:description: UVM testbench test
:files: /home/rrozak/antmicro/sv-tests/third_party/tests/easyUVM/top.sv
:incdirs: /home/rrozak/antmicro/sv-tests/third_party/tests/easyUVM
:tags: uvm
:timeout: 100
*/
